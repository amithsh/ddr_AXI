`include"common.sv"
`include "ddr_interface.sv"
`include"axi_interface.sv"
`include "ddr_cntrl.sv"
`include "dram.sv"
`include"axi_tx.sv"
`include"axi_gen.sv"
`include"axi_bfm.sv"
`include"AXI_slave_module.sv"
`include"axi_env.sv"
`include"axi_top.sv"
